`timescale 1ns/1ps
module routex_test();
   parameter STEP = 10;
   parameter Numports = 4;
   reg RST, CLK;

   reg [Numports-1:0][7:0][63:0]  D;
   reg [Numports-1:0]		  D_VALID;
   reg [Numports-1:0]		  Q_BP;
   
   wire [Numports-1:0][7:0][63:0] Q;
   
   reg [63:0]			  CNT;
   
   routex #(.PassThrough(4'b0)) uut (.RST(RST),
				     .CLK(CLK),
				     .D      (D),             // I [3:0][63:0]
				     .D_VALID(D_VALID),       // I [3:0]
				     .D_BP   (),              // O [3:0]
				     .Q       (Q),            // O [3:0][63:0]
				     .Q_VALID(),              // O [3:0]
				     .Q_BP   (Q_BP),          // I [3:0]
				     .Q_SOF   ());            // Not connected
   
   initial CLK <= 1;
   always #(STEP/2) CLK <= ~CLK;

   initial begin
      $shm_open();
      $shm_probe("ASM");

      RST <= 1;
      D <= 0;
      D_VALID <= 0;
      Q_BP <= 0;

      #(12.1*STEP)
      RST <= 0;
      
      #(1000*STEP)
      $finish;
   end // initial begin

   always @ (posedge CLK) begin
      if (RST) begin
	 CNT <= 0;
      end else begin 
	 CNT <= CNT + 1;
	 case (CNT)
	   101: begin
	      D[0][0] <= {8'h2, 56'h0};
	      D[0][1] <= {8'h2, 56'h0};
	      D[0][2] <= {8'h2, 56'h0};
	      D[0][3] <= {8'h1, 56'h1};
	      D[0][4] <= {8'h1, 56'h0};
	      D[0][5] <= {8'h1, 56'h0};
	      D[0][6] <= {8'h1, 56'h0};
	      D[0][7] <= 10;
	      
	      D[1][0] <= {8'h2, 56'h0};
	      D[1][1] <= {8'h2, 56'h0};
	      D[1][2] <= {8'h2, 56'h0};
	      D[1][3] <= {8'h1, 56'h1};
	      D[1][4] <= {8'h1, 56'h1};
	      D[1][5] <= {8'h1, 56'h1};
	      D[1][6] <= {8'h1, 56'h1};
	      D[1][7] <= 10;

	      D[2][0] <= {8'h2, 56'h1};
	      D[2][1] <= {8'h2, 56'h1};
	      D[2][2] <= {8'h2, 56'h1};
	      D[2][3] <= {8'h1, 56'h1};
	      D[2][4] <= {8'h1, 56'h1};
	      D[2][5] <= {8'h1, 56'h1};
	      D[2][6] <= {8'h1, 56'h1};
	      D[2][7] <= 10;

	      D[3][0] <= {8'h2, 56'h1};
	      D[3][1] <= {8'h2, 56'h1};
	      D[3][2] <= {8'h2, 56'h1};
	      D[3][3] <= {8'h1, 56'h1};
	      D[3][4] <= {8'h1, 56'h0};
	      D[3][5] <= {8'h1, 56'h0};
	      D[3][6] <= {8'h1, 56'h0};
	      D[3][7] <= 10;
	      
	      D_VALID[0] <= 1;
	      D_VALID[1] <= 1;
	      D_VALID[2] <= 1;
	      D_VALID[3] <= 1; end
	   101: begin
	      D[0][0] <= {8'h2, 56'h0};
	      D[0][1] <= {8'h2, 56'h0};
	      D[0][2] <= {8'h2, 56'h0};
	      D[0][3] <= {8'h1, 56'h1};
	      D[0][4] <= {8'h1, 56'h0};
	      D[0][5] <= {8'h1, 56'h0};
	      D[0][6] <= {8'h1, 56'h0};
	      D[0][7] <= 10;
	      
	      D[1][0] <= {8'h2, 56'h0};
	      D[1][1] <= {8'h2, 56'h0};
	      D[1][2] <= {8'h2, 56'h0};
	      D[1][3] <= {8'h1, 56'h1};
	      D[1][4] <= {8'h1, 56'h1};
	      D[1][5] <= {8'h1, 56'h1};
	      D[1][6] <= {8'h1, 56'h1};
	      D[1][7] <= 10;

	      D[2][0] <= {8'h2, 56'h1};
	      D[2][1] <= {8'h2, 56'h1};
	      D[2][2] <= {8'h2, 56'h1};
	      D[2][3] <= {8'h1, 56'h1};
	      D[2][4] <= {8'h1, 56'h1};
	      D[2][5] <= {8'h1, 56'h1};
	      D[2][6] <= {8'h1, 56'h1};
	      D[2][7] <= 10;

	      D[3][0] <= {8'h2, 56'h1};
	      D[3][1] <= {8'h2, 56'h1};
	      D[3][2] <= {8'h2, 56'h1};
	      D[3][3] <= {8'h1, 56'h1};
	      D[3][4] <= {8'h1, 56'h0};
	      D[3][5] <= {8'h1, 56'h0};
	      D[3][6] <= {8'h1, 56'h0};
	      D[3][7] <= 10;
	      
	      D_VALID[0] <= 1;
	      D_VALID[1] <= 1;
	      D_VALID[2] <= 1;
	      D_VALID[3] <= 1; end
	   102: begin
	      D[0][0] <= 64'h1;
	      D[0][1] <= 64'h2;
	      D[0][2] <= 64'h3;
	      D[0][3] <= 64'h4;
	      D[0][4] <= 64'h5;
	      D[0][5] <= 64'h6;
	      D[0][6] <= 64'h7;
	      D[0][7] <= 64'h8;

	      D[1][0] <= 64'h10;
	      D[1][1] <= 64'h20;
	      D[1][2] <= 64'h30;
	      D[1][3] <= 64'h40;
	      D[1][4] <= 64'h50;
	      D[1][5] <= 64'h60;
	      D[1][6] <= 64'h70;
	      D[1][7] <= 64'h80;
	      
	      D[2][0] <= 64'h100;
	      D[2][1] <= 64'h200;
	      D[2][2] <= 64'h300;
	      D[2][3] <= 64'h400;
	      D[2][4] <= 64'h500;
	      D[2][5] <= 64'h600;
	      D[2][6] <= 64'h700;
	      D[2][7] <= 64'h800;

	      D[3][0] <= 64'h1000;
	      D[3][1] <= 64'h2000;
	      D[3][2] <= 64'h3000;
	      D[3][3] <= 64'h4000;
	      D[3][4] <= 64'h5000;
	      D[3][5] <= 64'h6000;
	      D[3][6] <= 64'h7000;
	      D[3][7] <= 64'h8000; end
	   103: begin
	      D[0][0] <= 64'h9;
	      D[0][1] <= 64'h10;
	      
	      D[1][0] <= 64'h90;
	      D[1][1] <= 64'h100;

	      D[2][0] <= 64'h900;
	      D[2][1] <= 64'h1000;

	      D[3][0] <= 64'h9000;
	      D[3][1] <= 64'h10000; end
	   104: begin
	      D_VALID <= 0; end
	   201: begin
	      D[0][0] <= {8'h2, 56'h0};
	      D[0][1] <= {8'h2, 56'h3};
	      D[0][2] <= {8'h2, 56'h0};
	      D[0][3] <= {8'h2, 56'h0};
	      D[0][4] <= {8'h2, 56'h0};
	      D[0][5] <= {8'h2, 56'h0};
	      D[0][6] <= {8'h2, 56'h0};
	      D[0][7] <= {8'h2, 56'h3}; 
	      
	      D_VALID[0] <= 1;  end
	   202: begin
	      D[0][0] <= {8'h1, 56'h3};
	      D[0][1] <= {8'h1, 56'h0};
	      D[0][2] <= {8'h1, 56'h0};
	      D[0][3] <= {8'h1, 56'h0};
	      D[0][7] <= 32; end
	   203: begin
	      D[0][0] <= 64'h1;
	      D[0][1] <= 64'h2;
	      D[0][2] <= 64'h3;
	      D[0][3] <= 64'h4;
	      D[0][4] <= 64'h5;
	      D[0][5] <= 64'h6;
	      D[0][6] <= 64'h7;
	      D[0][7] <= 64'h8; end
	   204: begin 
	      D[0][0] <= 64'h9;
	      D[0][1] <= 64'h10;
	      D[0][2] <= 64'h11;
	      D[0][3] <= 64'h12;
	      D[0][4] <= 64'h13;
	      D[0][5] <= 64'h14;
	      D[0][6] <= 64'h15;
	      D[0][7] <= 64'h16; end
	   205: begin 
	      D[0][0] <= 64'h17;
	      D[0][1] <= 64'h18;
	      D[0][2] <= 64'h19;
	      D[0][3] <= 64'h20;
	      D[0][4] <= 64'h21;
	      D[0][5] <= 64'h22;
	      D[0][6] <= 64'h23;
	      D[0][7] <= 64'h24; end
	   206: begin 
	      D[0][0] <= 64'h25;
	      D[0][1] <= 64'h26;
	      D[0][2] <= 64'h27;
	      D[0][3] <= 64'h28;
	      D[0][4] <= 64'h29;
	      D[0][5] <= 64'h30;
	      D[0][6] <= 64'h31;
	      D[0][7] <= 64'h32; end
	   207: begin
	      D_VALID <= 0; end
	 endcase // case (CNT)
      end
   end // always @ (posedge CLK)
endmodule
