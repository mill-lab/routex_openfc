`timescale 1ns/1ps
module router_core_test();
   parameter STEP = 10;
   parameter Numports = 4;

   reg RST, CLK;

   reg [Numports-1:0][63:0] D;
   reg [Numports-1:0] 	    D_VALID;

   reg [63:0] 		    CNT;

   router_core #(.PassThrough(4'b0)) uut (.RST(RST),
					  .CLK(CLK),
					  .D(D),
					  .D_VALID(D_VALID),
					  .Q_BP(4'b0),
					  .D_BP(),
					  .COLLISION(),
					  .PT(),
					  .PT_VALID(),
					  .Q(),
					  .Q_VALID(),
					  .Q_SOF());

   initial CLK <= 1;
   always #(STEP/2) CLK <= ~CLK;

   initial begin
      $shm_open();
      $shm_probe("SA");

      RST <= 1;
      D <= 0;

      #(12.1*STEP)
      RST <= 0;

      #(100*STEP)
      $finish;
   end // initial begin

   always @ (posedge CLK) begin
      if (RST) begin
	 CNT <= 0;
      end else begin
	 CNT <= CNT + 1;
	 case (CNT)
	   1: begin
	      D[0] <= {8'h1, 56'h1};
	      D[1] <= {8'h1, 56'h1};
	      D_VALID[0] <= 1;
	      D_VALID[1] <= 1; end
	   2: begin
	      D[0] <= {8'h1, 56'h2};
	      D[1] <= {8'h1, 56'h2}; end
	   3: begin
	      D[0] <= 10;
	      D[1] <= 10; end
	   4: begin
	      D[0] <= 1;
	      D[1] <= 16*1;
	      D_VALID[1] <= 0; end
	   5: begin
	      D[0] <= 2;
	      D[1] <= {8'h1, 56'h1}; end
	   6: D[0] <= 3;
	   7: D[0] <= 4;
	   8: D[0] <= 5;
	   9: D[0] <= 6;
	   10: D[0] <= 7;
	   11: D[0] <= 8;
	   12: D[0] <= 9;
	   13: D[0] <= 10;
	   14: D_VALID[0] <= 0;
	   15:;
	   16:;
	   17:;
	   18:;
	   19:;
	   20:;
	   21:;
	   22:;
	   23: D_VALID[1] <= 1;
	   24: D[1] <= {8'h1, 56'h2};
	   25: D[1] <= 10;
	   26: D[1] <= 16*1;
	   27: D[1] <= 16*2;
	   28: D[1] <= 16*3;
	   29: D[1] <= 16*4;
	   30: D[1] <= 16*5;
	   31: D[1] <= 16*6;
	   32: D[1] <= 16*7;
	   33: D[1] <= 16*8;
	   34: D[1] <= 16*9;
	   35: D[1] <= 16*10;
	   36: D_VALID[1] <= 0;
	 endcase // case (CNT)
      end
   end // always @ (posedge CLK)
endmodule // router_core_test
