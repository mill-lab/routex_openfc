`timescale 1ns/1ps
`default_nettype none
module router_mux # (parameter NumPorts = 4, PortNo = 1) // n to 1 switch
   ( input wire CLK, RST,

     input wire [NumPorts-1:0][63:0] D,
     input wire [NumPorts-1:0][7:0]  DEST,
     input wire [NumPorts-1:0] 	     DEST_VALID, D_HDR_VALID, D_PLD_VALID,
     input wire [NumPorts-1:0] 	     D_SOF, D_EOF,
     output wire [NumPorts-1:0]      D_BP, COLLISION,

     output wire [63:0] 	     Q,
     output wire 		     Q_HDR_VALID, Q_PLD_VALID, Q_SOF, Q_EOF,
     input wire 		     Q_BP
     );

   genvar			     i;

   // - - - - - - - - - - - - - - - - - - - - 
   // SOF detection
   
   wire [NumPorts-1:0]           SOF_DETECT;

   generate
      for (i=0; i<NumPorts; i=i+1) begin : sof_detect_gen
         assign SOF_DETECT[i] = D_SOF[i] & (DEST[i] == PortNo);
      end
   endgenerate

   // - - - - - - - - - - - - - - - - - - - - 
   // Source switching on SOF_DETECT and corresponding EOF

   wire [NumPorts-1:0] SRC_PORTi;
   
   router_ch_sel # ( .NumCh(NumPorts) ) cs 
     ( .REQ(SOF_DETECT), .SEL(SRC_PORTi) );
   
   reg [NumPorts-1:0]  SRC_PORT;

   always @ (posedge CLK) begin
      if (RST) begin
         SRC_PORT <= 0;
      end else begin
         if (SRC_PORT==0) begin
            SRC_PORT <= SRC_PORTi;
         end else begin
            if (SRC_PORT & D_EOF) SRC_PORT <= 0;
         end
      end
   end

   // - - - - - - - - - - - - - - - - - - - -
   // Collision detection

   reg [NumPorts-1:0] CD;
   wire               EOF_DETECT = |(SRC_PORT & D_EOF);

   /*
   always @ (posedge CLK) begin
      if (RST) begin
         CD <= 0;
      end else begin
         CD <= (SRC_PORT==0) ? (SOF_DETECT & ~SRC_PORTi) :  // may be slow...
               (EOF_DETECT ? 0 :  // end of session
                CD | SOF_DETECT); // secondary collision 
      end
   end
    */

   reg [2:0]          EOF_CNT;
   wire               EOF_CNT_FULL = &EOF_CNT;
   
   always @ (posedge CLK) begin
      if (RST) begin
         CD <= 0;
         EOF_CNT <= 0;
      end else begin
         if (EOF_DETECT) EOF_CNT <= 1;
         else EOF_CNT <= (EOF_CNT != 0) ? EOF_CNT+1 : 0;

         if (CD==0) begin
            CD <= (SRC_PORT==0) ? (SOF_DETECT & ~SRC_PORTi) : 
                  (SOF_DETECT & ~SRC_PORT);
         end else begin
            CD <= EOF_CNT_FULL ? 0 : // end of session
                  CD | SOF_DETECT; // secondary collision
         end
      end

   end
    

   assign COLLISION = CD;
   
   // - - - - - - - - - - - - - - - - - - - - 
   // registered output

   wire [63:0] Qi_TMP;
   reg [63:0] Qi;
   reg        Q_HDR_VALIDi, Q_PLD_VALIDi, Q_SOFi, Q_EOFi;
   reg [NumPorts-1:0]  D_BPi;

   channel_mux # (.Width(64), .NumCh(NumPorts) ) dmux 
     ( .D(D), .SEL(SRC_PORT), .Q(Qi_TMP) );
   
   always @ (posedge CLK) begin
      Q_SOFi <= (SRC_PORT==0) & (|SOF_DETECT);
      Q_EOFi <= |(D_EOF & SRC_PORT);
      Q_HDR_VALIDi <= |(D_HDR_VALID & SRC_PORT);
      Q_PLD_VALIDi <= |(D_PLD_VALID & SRC_PORT);

      Qi <= Qi_TMP;
      D_BPi <= Q_BP ? SRC_PORT : 0;
   end
   
   assign Q     = Qi;
   assign Q_HDR_VALID = Q_HDR_VALIDi;
   assign Q_PLD_VALID = Q_PLD_VALIDi;
   assign Q_SOF = Q_SOFi;
   assign Q_EOF = Q_EOFi;
   assign D_BP  = D_BPi;
   
endmodule // router_mux
`default_nettype wire

// priprity circuit

module router_ch_sel # (parameter NumCh=8 )
   ( input wire [NumCh-1:0] REQ,
     output wire [NumCh-1:0] SEL );

   wire [NumCh-1:0][NumCh-1:0] TEMP;
   assign TEMP[0] = REQ[0] ? 1 : 0;
   
   generate
      genvar		       i;
      for (i=1; i<NumCh; i=i+1) begin : casex_gen
         assign TEMP[i] = (TEMP[i-1]!=0) ? TEMP[i-1] : (REQ[i] ? 1 << i : 0);
      end
   endgenerate

   assign SEL = TEMP[NumCh-1];
endmodule // channel_sel

// - - - - - - - - - - - - - - - - - - - - 
// Channel MUX with one-hot select signal

module channel_mux # ( parameter Width=64, NumCh=4 )
   ( input wire [NumCh-1:0][Width-1:0] D,
     input wire [NumCh-1:0]  SEL,
     output wire [Width-1:0] Q );
   
   wire [NumCh-1:0][Width-1:0] TEMP;
   
   assign TEMP[0] = SEL[0] ? D[0] : 0;

   generate
      genvar                   i;
      for (i=1; i<NumCh; i=i+1) begin : or_gen
         assign TEMP[i] = ( SEL[i] ? D[i] : 0) | TEMP[i-1];
      end
   endgenerate

   assign Q = TEMP[NumCh-1];
   
endmodule // channel_mux
